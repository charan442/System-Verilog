interface intf;
  logic d,q;
  logic clk,rst;
endinterface
