interface operation;
  logic a,b,c;
  logic sum, carry;
  
endinterface
