class transaction
  rand logic d;
  rand logic q;
  rand logic clk;
  rand logic rst;
  bit q;
endclass
