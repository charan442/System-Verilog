interface operation;
  logic clk;
  logic d;
  logic rst;
  bit q;
endinterface
