class transaction;
  randc logic d;
  bit q;
endclass
